`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:08:05 01/14/2015 
// Design Name: 
// Module Name:    segment_translater 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module segment_translater(
input CLK
//	output [7:0] digitOneTranslated,
//	output [7:0] digitTwoTranslated,
//	output [7:0] digitThreeTranslated,
//	output [7:0] digitFourTranslated
    );


endmodule
